`timescale 1ns/1ps
`default_nettype none

module top_level (
    input wire a,
    input wire [] b,
    output logic c,
);
    
endmodule
`default_nettype wire ;